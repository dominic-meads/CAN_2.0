////////////////////////////////////////////////////////////////////////////////
// Copyright (C) 1999-2008 Easics NV.
// This source file may be used and distributed without restriction
// provided that this copyright statement is not removed from the file
// and that any derivative work contains the original copyright notice
// and the associated disclaimer.
//
// THIS SOURCE FILE IS PROVIDED "AS IS" AND WITHOUT ANY EXPRESS
// OR IMPLIED WARRANTIES, INCLUDING, WITHOUT LIMITATION, THE IMPLIED
// WARRANTIES OF MERCHANTIBILITY AND FITNESS FOR A PARTICULAR PURPOSE.
//
// Purpose : synthesizable CRC function
//   * polynomial: x^15 + x^14 + x^10 + x^8 + x^7 + x^4 + x^3 + x^1 + 1
//   * data width: 83
//
// Info : tools@easics.be
//        http://www.easics.com
////////////////////////////////////////////////////////////////////////////////
`timescale 1 ns / 1 ps
module CRC15_D83(
 // input clk,
 // input rst_n,
  input reg [82:0] din,
  output [14:0] o_crc
);
  
  reg [14:0] r_seed = 15'hFFFF;  // Must be seeded with all 1's 
  reg [14:0] r_crc;

  // polynomial: x^15 + x^14 + x^10 + x^8 + x^7 + x^4 + x^3 + x^1 + 1
  // data width: 83
  // convention: the first serial bit is D[82]
  function [14:0] nextCRC15_D83;

    input [82:0] Data;
    input [14:0] crc;
    reg [82:0] d;
    reg [14:0] c;
    reg [14:0] newcrc;
  begin
    d = Data;
    c = crc;

    newcrc[0] = d[82] ^ d[79] ^ d[77] ^ d[76] ^ d[75] ^ d[73] ^ d[72] ^ d[70] ^ d[66] ^ d[65] ^ d[64] ^ d[63] ^ d[62] ^ d[61] ^ d[60] ^ d[59] ^ d[58] ^ d[53] ^ d[52] ^ d[50] ^ d[47] ^ d[46] ^ d[45] ^ d[44] ^ d[40] ^ d[37] ^ d[36] ^ d[35] ^ d[34] ^ d[33] ^ d[27] ^ d[26] ^ d[22] ^ d[21] ^ d[19] ^ d[18] ^ d[17] ^ d[16] ^ d[12] ^ d[11] ^ d[10] ^ d[9] ^ d[7] ^ d[6] ^ d[4] ^ d[3] ^ d[2] ^ d[1] ^ d[0] ^ c[2] ^ c[4] ^ c[5] ^ c[7] ^ c[8] ^ c[9] ^ c[11] ^ c[14];
    newcrc[1] = d[82] ^ d[80] ^ d[79] ^ d[78] ^ d[75] ^ d[74] ^ d[72] ^ d[71] ^ d[70] ^ d[67] ^ d[58] ^ d[54] ^ d[52] ^ d[51] ^ d[50] ^ d[48] ^ d[44] ^ d[41] ^ d[40] ^ d[38] ^ d[33] ^ d[28] ^ d[26] ^ d[23] ^ d[21] ^ d[20] ^ d[16] ^ d[13] ^ d[9] ^ d[8] ^ d[6] ^ d[5] ^ d[0] ^ c[2] ^ c[3] ^ c[4] ^ c[6] ^ c[7] ^ c[10] ^ c[11] ^ c[12] ^ c[14];
    newcrc[2] = d[81] ^ d[80] ^ d[79] ^ d[76] ^ d[75] ^ d[73] ^ d[72] ^ d[71] ^ d[68] ^ d[59] ^ d[55] ^ d[53] ^ d[52] ^ d[51] ^ d[49] ^ d[45] ^ d[42] ^ d[41] ^ d[39] ^ d[34] ^ d[29] ^ d[27] ^ d[24] ^ d[22] ^ d[21] ^ d[17] ^ d[14] ^ d[10] ^ d[9] ^ d[7] ^ d[6] ^ d[1] ^ c[0] ^ c[3] ^ c[4] ^ c[5] ^ c[7] ^ c[8] ^ c[11] ^ c[12] ^ c[13];
    newcrc[3] = d[81] ^ d[80] ^ d[79] ^ d[75] ^ d[74] ^ d[70] ^ d[69] ^ d[66] ^ d[65] ^ d[64] ^ d[63] ^ d[62] ^ d[61] ^ d[59] ^ d[58] ^ d[56] ^ d[54] ^ d[47] ^ d[45] ^ d[44] ^ d[43] ^ d[42] ^ d[37] ^ d[36] ^ d[34] ^ d[33] ^ d[30] ^ d[28] ^ d[27] ^ d[26] ^ d[25] ^ d[23] ^ d[21] ^ d[19] ^ d[17] ^ d[16] ^ d[15] ^ d[12] ^ d[9] ^ d[8] ^ d[6] ^ d[4] ^ d[3] ^ d[1] ^ d[0] ^ c[1] ^ c[2] ^ c[6] ^ c[7] ^ c[11] ^ c[12] ^ c[13];
    newcrc[4] = d[81] ^ d[80] ^ d[79] ^ d[77] ^ d[73] ^ d[72] ^ d[71] ^ d[67] ^ d[61] ^ d[58] ^ d[57] ^ d[55] ^ d[53] ^ d[52] ^ d[50] ^ d[48] ^ d[47] ^ d[43] ^ d[40] ^ d[38] ^ d[36] ^ d[33] ^ d[31] ^ d[29] ^ d[28] ^ d[24] ^ d[21] ^ d[20] ^ d[19] ^ d[13] ^ d[12] ^ d[11] ^ d[6] ^ d[5] ^ d[3] ^ d[0] ^ c[3] ^ c[4] ^ c[5] ^ c[9] ^ c[11] ^ c[12] ^ c[13];
    newcrc[5] = d[82] ^ d[81] ^ d[80] ^ d[78] ^ d[74] ^ d[73] ^ d[72] ^ d[68] ^ d[62] ^ d[59] ^ d[58] ^ d[56] ^ d[54] ^ d[53] ^ d[51] ^ d[49] ^ d[48] ^ d[44] ^ d[41] ^ d[39] ^ d[37] ^ d[34] ^ d[32] ^ d[30] ^ d[29] ^ d[25] ^ d[22] ^ d[21] ^ d[20] ^ d[14] ^ d[13] ^ d[12] ^ d[7] ^ d[6] ^ d[4] ^ d[1] ^ c[0] ^ c[4] ^ c[5] ^ c[6] ^ c[10] ^ c[12] ^ c[13] ^ c[14];
    newcrc[6] = d[82] ^ d[81] ^ d[79] ^ d[75] ^ d[74] ^ d[73] ^ d[69] ^ d[63] ^ d[60] ^ d[59] ^ d[57] ^ d[55] ^ d[54] ^ d[52] ^ d[50] ^ d[49] ^ d[45] ^ d[42] ^ d[40] ^ d[38] ^ d[35] ^ d[33] ^ d[31] ^ d[30] ^ d[26] ^ d[23] ^ d[22] ^ d[21] ^ d[15] ^ d[14] ^ d[13] ^ d[8] ^ d[7] ^ d[5] ^ d[2] ^ c[1] ^ c[5] ^ c[6] ^ c[7] ^ c[11] ^ c[13] ^ c[14];
    newcrc[7] = d[80] ^ d[79] ^ d[77] ^ d[74] ^ d[73] ^ d[72] ^ d[66] ^ d[65] ^ d[63] ^ d[62] ^ d[59] ^ d[56] ^ d[55] ^ d[52] ^ d[51] ^ d[47] ^ d[45] ^ d[44] ^ d[43] ^ d[41] ^ d[40] ^ d[39] ^ d[37] ^ d[35] ^ d[33] ^ d[32] ^ d[31] ^ d[26] ^ d[24] ^ d[23] ^ d[21] ^ d[19] ^ d[18] ^ d[17] ^ d[15] ^ d[14] ^ d[12] ^ d[11] ^ d[10] ^ d[8] ^ d[7] ^ d[4] ^ d[2] ^ d[1] ^ d[0] ^ c[4] ^ c[5] ^ c[6] ^ c[9] ^ c[11] ^ c[12];
    newcrc[8] = d[82] ^ d[81] ^ d[80] ^ d[79] ^ d[78] ^ d[77] ^ d[76] ^ d[74] ^ d[72] ^ d[70] ^ d[67] ^ d[65] ^ d[62] ^ d[61] ^ d[59] ^ d[58] ^ d[57] ^ d[56] ^ d[50] ^ d[48] ^ d[47] ^ d[42] ^ d[41] ^ d[38] ^ d[37] ^ d[35] ^ d[32] ^ d[26] ^ d[25] ^ d[24] ^ d[21] ^ d[20] ^ d[17] ^ d[15] ^ d[13] ^ d[10] ^ d[8] ^ d[7] ^ d[6] ^ d[5] ^ d[4] ^ d[0] ^ c[2] ^ c[4] ^ c[6] ^ c[8] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[14];
    newcrc[9] = d[82] ^ d[81] ^ d[80] ^ d[79] ^ d[78] ^ d[77] ^ d[75] ^ d[73] ^ d[71] ^ d[68] ^ d[66] ^ d[63] ^ d[62] ^ d[60] ^ d[59] ^ d[58] ^ d[57] ^ d[51] ^ d[49] ^ d[48] ^ d[43] ^ d[42] ^ d[39] ^ d[38] ^ d[36] ^ d[33] ^ d[27] ^ d[26] ^ d[25] ^ d[22] ^ d[21] ^ d[18] ^ d[16] ^ d[14] ^ d[11] ^ d[9] ^ d[8] ^ d[7] ^ d[6] ^ d[5] ^ d[1] ^ c[0] ^ c[3] ^ c[5] ^ c[7] ^ c[9] ^ c[10] ^ c[11] ^ c[12] ^ c[13] ^ c[14];
    newcrc[10] = d[81] ^ d[80] ^ d[78] ^ d[77] ^ d[75] ^ d[74] ^ d[73] ^ d[70] ^ d[69] ^ d[67] ^ d[66] ^ d[65] ^ d[62] ^ d[53] ^ d[49] ^ d[47] ^ d[46] ^ d[45] ^ d[43] ^ d[39] ^ d[36] ^ d[35] ^ d[33] ^ d[28] ^ d[23] ^ d[21] ^ d[18] ^ d[16] ^ d[15] ^ d[11] ^ d[8] ^ d[4] ^ d[3] ^ d[1] ^ d[0] ^ c[1] ^ c[2] ^ c[5] ^ c[6] ^ c[7] ^ c[9] ^ c[10] ^ c[12] ^ c[13];
    newcrc[11] = d[82] ^ d[81] ^ d[79] ^ d[78] ^ d[76] ^ d[75] ^ d[74] ^ d[71] ^ d[70] ^ d[68] ^ d[67] ^ d[66] ^ d[63] ^ d[54] ^ d[50] ^ d[48] ^ d[47] ^ d[46] ^ d[44] ^ d[40] ^ d[37] ^ d[36] ^ d[34] ^ d[29] ^ d[24] ^ d[22] ^ d[19] ^ d[17] ^ d[16] ^ d[12] ^ d[9] ^ d[5] ^ d[4] ^ d[2] ^ d[1] ^ c[0] ^ c[2] ^ c[3] ^ c[6] ^ c[7] ^ c[8] ^ c[10] ^ c[11] ^ c[13] ^ c[14];
    newcrc[12] = d[82] ^ d[80] ^ d[79] ^ d[77] ^ d[76] ^ d[75] ^ d[72] ^ d[71] ^ d[69] ^ d[68] ^ d[67] ^ d[64] ^ d[55] ^ d[51] ^ d[49] ^ d[48] ^ d[47] ^ d[45] ^ d[41] ^ d[38] ^ d[37] ^ d[35] ^ d[30] ^ d[25] ^ d[23] ^ d[20] ^ d[18] ^ d[17] ^ d[13] ^ d[10] ^ d[6] ^ d[5] ^ d[3] ^ d[2] ^ c[0] ^ c[1] ^ c[3] ^ c[4] ^ c[7] ^ c[8] ^ c[9] ^ c[11] ^ c[12] ^ c[14];
    newcrc[13] = d[81] ^ d[80] ^ d[78] ^ d[77] ^ d[76] ^ d[73] ^ d[72] ^ d[70] ^ d[69] ^ d[68] ^ d[65] ^ d[56] ^ d[52] ^ d[50] ^ d[49] ^ d[48] ^ d[46] ^ d[42] ^ d[39] ^ d[38] ^ d[36] ^ d[31] ^ d[26] ^ d[24] ^ d[21] ^ d[19] ^ d[18] ^ d[14] ^ d[11] ^ d[7] ^ d[6] ^ d[4] ^ d[3] ^ c[0] ^ c[1] ^ c[2] ^ c[4] ^ c[5] ^ c[8] ^ c[9] ^ c[10] ^ c[12] ^ c[13];
    newcrc[14] = d[81] ^ d[78] ^ d[76] ^ d[75] ^ d[74] ^ d[72] ^ d[71] ^ d[69] ^ d[65] ^ d[64] ^ d[63] ^ d[62] ^ d[61] ^ d[60] ^ d[59] ^ d[58] ^ d[57] ^ d[52] ^ d[51] ^ d[49] ^ d[46] ^ d[45] ^ d[44] ^ d[43] ^ d[39] ^ d[36] ^ d[35] ^ d[34] ^ d[33] ^ d[32] ^ d[26] ^ d[25] ^ d[21] ^ d[20] ^ d[18] ^ d[17] ^ d[16] ^ d[15] ^ d[11] ^ d[10] ^ d[9] ^ d[8] ^ d[6] ^ d[5] ^ d[3] ^ d[2] ^ d[1] ^ d[0] ^ c[1] ^ c[3] ^ c[4] ^ c[6] ^ c[7] ^ c[8] ^ c[10] ^ c[13];
    nextCRC15_D83 = newcrc;
  end
  endfunction
  
  always @ (*)
    begin 
      if (!rst_n)
        begin
          r_seed = 15'hFFFF;
          r_crc = 15'h0000;
        end 
      else 
        begin
          o_crc = nextCRC15_D83(din, r_seed);
        end
      
endmodule
